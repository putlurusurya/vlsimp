magic
tech min2
timestamp 1606752020
<< nwell >>
rect -13 24 26 69
<< ntransistor >>
rect 1 1 3 6
rect 10 1 12 6
<< ptransistor >>
rect 1 47 3 57
rect 10 47 12 57
<< ndiffusion >>
rect -4 5 1 6
rect 0 1 1 5
rect 3 2 4 6
rect 9 2 10 6
rect 3 1 10 2
rect 12 5 17 6
rect 12 1 13 5
<< pdiffusion >>
rect 0 53 1 57
rect -4 52 1 53
rect 0 48 1 52
rect -4 47 1 48
rect 3 47 10 57
rect 12 56 17 57
rect 12 52 13 56
rect 12 51 17 52
rect 12 47 13 51
<< ndcontact >>
rect -4 1 0 5
rect 4 2 9 6
rect 13 1 17 5
<< pdcontact >>
rect -4 53 0 57
rect -4 48 0 52
rect 13 52 17 56
rect 13 47 17 51
<< psubstratepcontact >>
rect -11 -7 -7 -3
rect 5 -7 9 -3
rect 20 -7 24 -3
<< nsubstratencontact >>
rect -10 61 -6 65
rect 5 61 9 65
rect 19 61 23 65
<< polysilicon >>
rect 1 57 3 59
rect 10 57 12 59
rect 1 6 3 47
rect 10 6 12 47
rect 1 -1 3 1
rect 10 -1 12 1
<< polycontact >>
rect -3 34 1 38
rect 6 28 10 32
<< metal1 >>
rect -11 61 -10 65
rect -6 61 5 65
rect 9 61 19 65
rect 23 61 24 65
rect -11 59 24 61
rect -4 57 0 59
rect -4 52 0 53
rect 13 51 17 52
rect -4 34 -3 38
rect 5 28 6 32
rect 13 19 17 47
rect 5 15 24 19
rect 5 6 8 15
rect -4 -1 0 1
rect 13 -1 17 1
rect -11 -3 24 -1
rect -7 -7 5 -3
rect 9 -7 20 -3
<< labels >>
rlabel metal1 2 -4 2 -4 1 Gnd
rlabel metal1 24 15 24 19 7 out
rlabel metal1 2 63 2 63 5 vdd
rlabel polycontact -1 36 -1 36 1 a
rlabel polycontact 8 30 8 30 1 b
<< end >>
