magic
tech min2
timestamp 1606801835
<< nwell >>
rect -12 24 22 68
<< ntransistor >>
rect 1 3 3 8
rect 6 3 8 8
<< ptransistor >>
rect 1 45 3 55
rect 6 45 8 55
<< ndiffusion >>
rect -4 7 1 8
rect 0 3 1 7
rect 3 3 6 8
rect 8 4 9 8
rect 8 3 13 4
<< pdiffusion >>
rect -4 50 1 55
rect 0 46 1 50
rect -4 45 1 46
rect 3 45 6 55
rect 8 53 13 55
rect 8 49 9 53
rect 8 45 13 49
<< ndcontact >>
rect -4 3 0 7
rect 9 4 13 8
<< pdcontact >>
rect -4 46 0 50
rect 9 49 13 53
<< psubstratepcontact >>
rect -11 -7 -7 -3
rect 10 -7 14 -3
<< nsubstratencontact >>
rect -9 61 -5 65
rect 10 61 14 65
<< polysilicon >>
rect 1 57 8 59
rect 1 55 3 57
rect 6 55 8 57
rect 1 8 3 45
rect 6 8 8 45
rect 1 1 3 3
rect 6 1 8 3
rect 1 -1 8 1
<< polycontact >>
rect -3 16 1 20
<< metal1 >>
rect -11 61 -9 65
rect -5 61 10 65
rect 14 61 21 65
rect -11 59 21 61
rect -4 50 0 59
rect 9 53 13 54
rect 9 28 13 49
rect 9 24 21 28
rect -4 16 -3 20
rect 9 8 13 24
rect -4 -1 0 3
rect -11 -3 21 -1
rect -7 -7 10 -3
rect 14 -7 21 -3
<< labels >>
rlabel polycontact -1 18 -1 18 1 a
rlabel metal1 2 -4 2 -4 1 Gnd
rlabel metal1 2 63 2 63 5 vdd
rlabel metal1 21 24 21 28 7 out
<< end >>
