* SPICE3 file created from and.ext - technology: min2

.option scale=0.1u

M1000 a_n17_1# b vdd vdd pfet w=10 l=2
+  ad=70 pd=34 as=120 ps=64
M1001 vdd a a_n17_1# vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_8_47# a_n17_1# vdd vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1003 a_13_47# a_n17_1# a_8_47# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1004 a_18_47# a_n17_1# a_13_47# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1005 out a_n17_1# a_18_47# vdd pfet w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1006 a_n10_1# b a_n17_1# Gnd nfet w=5 l=2
+  ad=35 pd=24 as=25 ps=20
M1007 Gnd a a_n10_1# Gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1008 a_8_1# a_n17_1# Gnd Gnd nfet w=5 l=2
+  ad=15 pd=16 as=0 ps=0
M1009 a_13_1# a_n17_1# a_8_1# Gnd nfet w=5 l=2
+  ad=15 pd=16 as=0 ps=0
M1010 a_18_1# a_n17_1# a_13_1# Gnd nfet w=5 l=2
+  ad=15 pd=16 as=0 ps=0
M1011 out a_n17_1# a_18_1# Gnd nfet w=5 l=2
+  ad=30 pd=22 as=0 ps=0
C0 vdd b 0.18482fF
C1 vdd a 0.18482fF
C2 b a 0.16295fF
C3 vdd a_n17_1# 1.14232fF
C4 b a_n17_1# 0.07186fF
C5 a a_n17_1# 0.22979fF
C6 vdd out 0.16569fF
C7 vdd Gnd 0.00202fF


.include NMOS-180nm.lib
.include PMOS-180nm.lib


v_dd vdd Gnd 1.8
v_d a Gnd pulse( 1.8 0 0 1ns 1ns 50ns 100ns)

v1 b Gnd pulse(1.8 0 0 1ns 1ns 100ns 200ns)

.control
	tran 0.1ns 200ns
	
	plot tran1.a tran1.b tran1.out
	
	meas tran risetime  trig out val=0.18 RISE=1 TARG out val=1.62 RISE=1

	meas tran falltime  trig out val=1.62  FALL=1 TARG out val=0.18 FALL=1
	
	meas tran tplh trig a val=0.9 RISE=2 TARG out val=0.9 RISE=1
	
	meas tran tphl trig a val=0.9 FALL=1 TARG out val=0.9 FALL=1
	
	let x= -tran1.v_dd#branch
        
        plot vdd*x	   
	    
.endc

