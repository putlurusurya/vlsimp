* SPICE3 file created from nand.ext - technology: min2

.option scale=0.1u

.include NMOS-180nm.lib
.include PMOS-180nm.lib
M1000 out a vdd vdd pfet w=10 l=2
+  ad=70 pd=34 as=100 ps=60
M1001 vdd b out vdd pfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_3_1# a Gnd Gnd nfet w=5 l=2
+  ad=35 pd=24 as=25 ps=20
M1003 out b a_3_1# Gnd nfet w=5 l=2
+  ad=25 pd=20 as=0 ps=0
C0 vdd a 0.18482fF
C1 vdd b 0.18482fF
C2 vdd out 0.34494fF
C3 a b 0.6295fF
C4 b out 0.07186fF

v1 vdd Gnd 1.8
vin1 a Gnd pulse( 1.8 0 0 1n 1n 20n 50n)
vin2 b Gnd pulse( 1.8 0 0 1n 1n 40n 80n)

.tran 0.1n 200n

.control
	tran 0.1ns 200ns
	
	plot tran1.a tran1.b tran1.out
	
	meas tran risetime  trig out val=0.18 RISE=1 TARG out val=1.62 RISE=1

	meas tran falltime  trig out val=1.62  FALL=1 TARG out val=0.18 FALL=1
	
	meas tran tplh trig a val=0.9 FALL=1 TARG out val=0.9 RISE=1
	
	meas tran tphl trig b val=0.9 RISE=1 TARG out val=0.9 FALL=1
	
	let x= -tran1.v1#branch
        
        plot vdd*x	   
	    
.endc
