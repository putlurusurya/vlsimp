* SPICE3 file created from inverter.ext - technology: min2

.option scale=0.1u

.include NMOS-180nm.lib
.include PMOS-180nm.lib
M1000 out a vdd vdd pfet w=10 l=2
+  ad=50 pd=30 as=50 ps=30
M1001 out a Gnd Gnd nfet w=5 l=2
+  ad=25 pd=20 as=25 ps=20
C0 a out 0.05498fF
C1 vdd a 0.18482fF
C2 vdd out 0.25929fF



v1 vdd Gnd 1.8
vin1 a Gnd pulse(0 1.8 0 1n 1n 30n 60n)

.tran 0.1n 200n

.control
run

meas tran risetime  trig out val=0.18 RISE=1 TARG out val=1.62 RISE=1

meas tran falltime  trig out val=1.62  FALL=1 TARG out val=0.18 FALL=1

meas tran tphl trig a val=0.9  RISE=1 TARG out val=0.9 FALL=1

meas tran tplh trig a val=0.9  FALL=1 TARG out val=0.9 RISE=1

plot V(a)  V(out)

let x= -tran1.v1#branch
        
        plot vdd*x
.endc
