magic
tech min2
timestamp 1606884912
<< nwell >>
rect -52 24 28 69
<< ntransistor >>
rect -39 1 -37 6
rect -34 1 -32 6
rect -29 1 -27 6
rect -24 1 -22 6
rect -6 1 -4 6
rect 2 1 4 6
rect 11 1 13 6
<< ptransistor >>
rect -39 47 -37 57
rect -34 47 -32 57
rect -29 47 -27 57
rect -24 47 -22 57
rect -6 47 -4 57
rect 2 47 4 57
rect 11 47 13 57
<< ndiffusion >>
rect -41 2 -39 6
rect -45 1 -39 2
rect -37 1 -34 6
rect -32 1 -29 6
rect -27 1 -24 6
rect -22 5 -16 6
rect -22 1 -20 5
rect -8 2 -6 6
rect -12 1 -6 2
rect -4 5 2 6
rect -4 1 -3 5
rect 1 1 2 5
rect 4 1 11 6
rect 13 2 14 6
rect 13 1 18 2
<< pdiffusion >>
rect -45 56 -39 57
rect -41 52 -39 56
rect -45 51 -39 52
rect -41 47 -39 51
rect -37 47 -34 57
rect -32 47 -29 57
rect -27 47 -24 57
rect -22 53 -20 57
rect -22 52 -16 53
rect -22 48 -20 52
rect -22 47 -16 48
rect -12 56 -6 57
rect -8 52 -6 56
rect -12 51 -6 52
rect -8 47 -6 51
rect -4 52 2 57
rect -4 48 -3 52
rect 1 48 2 52
rect -4 47 2 48
rect 4 55 11 57
rect 4 51 5 55
rect 10 51 11 55
rect 4 47 11 51
rect 13 52 18 57
rect 13 48 14 52
rect 13 47 18 48
<< ndcontact >>
rect -45 2 -41 6
rect -20 1 -16 5
rect -12 2 -8 6
rect -3 1 1 5
rect 14 2 18 6
<< pdcontact >>
rect -45 52 -41 56
rect -45 47 -41 51
rect -20 53 -16 57
rect -20 48 -16 52
rect -12 52 -8 56
rect -12 47 -8 51
rect -3 48 1 52
rect 5 51 10 55
rect 14 48 18 52
<< psubstratepcontact >>
rect -49 -7 -45 -3
rect 6 -7 10 -3
rect 21 -7 25 -3
<< nsubstratencontact >>
rect -49 61 -45 65
rect 6 61 10 65
rect 21 61 25 65
<< polysilicon >>
rect -39 57 -37 59
rect -34 57 -32 59
rect -29 57 -27 59
rect -24 57 -22 59
rect -6 57 -4 59
rect 2 57 4 59
rect 11 57 13 59
rect -39 45 -37 47
rect -34 45 -32 47
rect -29 45 -27 47
rect -24 45 -22 47
rect -39 41 -22 45
rect -39 14 -37 41
rect -34 14 -32 41
rect -29 14 -27 41
rect -24 28 -22 41
rect -6 31 -4 47
rect -24 24 -23 28
rect -6 27 -5 31
rect -24 14 -22 24
rect -39 10 -22 14
rect -39 6 -37 10
rect -34 6 -32 10
rect -29 6 -27 10
rect -24 6 -22 10
rect -6 6 -4 27
rect 2 20 4 47
rect 3 16 4 20
rect 2 6 4 16
rect 11 6 13 47
rect -39 -1 -37 1
rect -34 -1 -32 1
rect -29 -1 -27 1
rect -24 -1 -22 1
rect -6 -1 -4 1
rect 2 -1 4 1
rect 11 -1 13 1
<< polycontact >>
rect -23 24 -19 28
rect -5 27 -1 31
rect -1 16 3 20
rect 7 12 11 16
<< metal1 >>
rect -45 61 6 65
rect 10 61 21 65
rect -49 59 25 61
rect -20 57 -16 59
rect -45 51 -41 52
rect -20 52 -16 53
rect -12 51 -8 52
rect -45 6 -41 47
rect -3 52 1 59
rect 6 55 9 56
rect 14 52 18 59
rect -12 28 -8 47
rect 6 31 9 51
rect -19 24 -8 28
rect -1 27 18 31
rect -12 6 -8 24
rect -2 16 -1 20
rect 6 12 7 16
rect 14 6 18 27
rect -20 -1 -16 1
rect -3 -1 1 1
rect -49 -3 25 -1
rect -45 -7 6 -3
rect 10 -7 21 -3
<< labels >>
rlabel polycontact 9 14 9 14 1 b
rlabel metal1 3 -4 3 -4 1 Gnd
rlabel metal1 3 63 3 63 5 vdd
rlabel polycontact 1 18 1 18 1 a
rlabel metal1 -43 26 -43 26 1 out
<< end >>
