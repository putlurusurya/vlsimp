magic
tech min2
timestamp 1606899548
<< nwell >>
rect -26 31 91 75
<< ntransistor >>
rect -14 18 -12 25
rect -4 18 -2 25
rect 13 18 15 25
rect 21 18 23 25
rect 32 18 34 23
rect 41 18 43 25
rect 49 18 51 25
rect 57 18 59 25
rect 69 18 71 23
rect 78 18 80 25
<< ptransistor >>
rect -14 39 -12 53
rect -4 39 -2 53
rect 13 39 15 53
rect 21 39 23 53
rect 32 39 34 48
rect 41 39 43 53
rect 49 39 51 53
rect 57 39 59 53
rect 69 39 71 48
rect 78 39 80 53
<< ndiffusion >>
rect -20 24 -14 25
rect -16 19 -14 24
rect -20 18 -14 19
rect -12 24 -4 25
rect -12 19 -10 24
rect -6 19 -4 24
rect -12 18 -4 19
rect -2 24 4 25
rect -2 19 0 24
rect -2 18 4 19
rect 8 24 13 25
rect 12 19 13 24
rect 8 18 13 19
rect 15 19 16 25
rect 20 19 21 25
rect 15 18 21 19
rect 23 23 29 25
rect 36 23 41 25
rect 23 19 25 23
rect 29 19 32 23
rect 23 18 32 19
rect 34 18 36 23
rect 40 18 41 23
rect 43 19 44 25
rect 48 19 49 25
rect 43 18 49 19
rect 51 19 52 25
rect 56 19 57 25
rect 51 18 57 19
rect 59 23 66 25
rect 73 23 78 25
rect 59 19 62 23
rect 66 19 69 23
rect 59 18 69 19
rect 71 18 73 23
rect 77 18 78 23
rect 80 20 81 25
rect 80 18 85 20
<< pdiffusion >>
rect -20 52 -14 53
rect -16 47 -14 52
rect -20 44 -14 47
rect -16 39 -14 44
rect -12 52 -4 53
rect -12 47 -10 52
rect -6 47 -4 52
rect -12 44 -4 47
rect -12 39 -10 44
rect -6 39 -4 44
rect -2 52 4 53
rect -2 47 0 52
rect -2 44 4 47
rect -2 39 0 44
rect 8 52 13 53
rect 12 47 13 52
rect 8 44 13 47
rect 12 39 13 44
rect 15 52 21 53
rect 15 48 16 52
rect 20 48 21 52
rect 15 43 21 48
rect 15 39 16 43
rect 20 39 21 43
rect 23 52 29 53
rect 23 48 25 52
rect 40 49 41 53
rect 36 48 41 49
rect 23 47 32 48
rect 23 41 25 47
rect 29 41 32 47
rect 23 39 32 41
rect 34 44 41 48
rect 34 40 36 44
rect 40 40 41 44
rect 34 39 41 40
rect 43 52 49 53
rect 43 48 44 52
rect 48 48 49 52
rect 43 43 49 48
rect 43 39 44 43
rect 48 39 49 43
rect 51 52 57 53
rect 51 48 52 52
rect 56 48 57 52
rect 51 43 57 48
rect 51 39 52 43
rect 56 39 57 43
rect 59 52 66 53
rect 59 48 62 52
rect 77 49 78 53
rect 73 48 78 49
rect 59 47 69 48
rect 59 41 62 47
rect 66 41 69 47
rect 59 39 69 41
rect 71 44 78 48
rect 71 40 73 44
rect 77 40 78 44
rect 71 39 78 40
rect 80 52 85 53
rect 80 48 81 52
rect 80 43 85 48
rect 80 39 81 43
<< ndcontact >>
rect -20 19 -16 24
rect -10 19 -6 24
rect 0 19 4 24
rect 8 19 12 24
rect 16 19 20 25
rect 25 19 29 23
rect 36 18 40 23
rect 44 19 48 25
rect 52 19 56 25
rect 62 19 66 23
rect 73 18 77 23
rect 81 20 85 25
<< pdcontact >>
rect -20 47 -16 52
rect -20 39 -16 44
rect -10 47 -6 52
rect -10 39 -6 44
rect 0 47 4 52
rect 0 39 4 44
rect 8 47 12 52
rect 8 39 12 44
rect 16 48 20 52
rect 16 39 20 43
rect 25 48 29 52
rect 36 49 40 53
rect 25 41 29 47
rect 36 40 40 44
rect 44 48 48 52
rect 44 39 48 43
rect 52 48 56 52
rect 52 39 56 43
rect 62 48 66 52
rect 73 49 77 53
rect 62 41 66 47
rect 73 40 77 44
rect 81 48 85 52
rect 81 39 85 43
<< nsubstratendiff >>
rect 25 68 29 72
rect 47 68 53 72
rect 63 68 67 72
<< psubstratepcontact >>
rect 1 0 5 4
rect 17 0 21 4
rect 36 0 40 4
rect 57 0 61 4
rect 79 0 83 4
<< nsubstratencontact >>
rect 3 68 7 72
rect 17 68 21 72
rect 29 68 35 72
rect 53 68 57 72
rect 67 68 72 72
rect 81 68 85 72
<< polysilicon >>
rect -16 62 7 64
rect -16 60 -12 62
rect -14 53 -12 60
rect -4 53 -2 55
rect -14 37 -12 39
rect -4 33 -2 39
rect -14 31 -2 33
rect -14 25 -12 31
rect -4 25 -2 27
rect -14 13 -12 18
rect -4 12 -2 18
rect 5 12 7 62
rect 24 64 51 66
rect 12 54 15 56
rect 13 53 15 54
rect 21 53 23 61
rect 31 59 43 61
rect 41 53 43 59
rect 49 53 51 64
rect 68 59 80 61
rect 57 53 59 55
rect 78 53 80 59
rect 32 48 34 50
rect 69 48 71 50
rect 13 34 15 39
rect 21 37 23 39
rect 32 35 34 39
rect 13 32 23 34
rect 13 25 15 27
rect 21 25 23 32
rect 32 23 34 30
rect 41 25 43 39
rect 49 37 51 39
rect 57 34 59 39
rect 49 32 59 34
rect 69 35 71 39
rect 49 25 51 32
rect 57 25 59 27
rect 69 23 71 30
rect 78 25 80 39
rect -4 10 7 12
rect 13 11 15 18
rect 21 13 23 18
rect 32 16 34 18
rect 41 16 43 18
rect 49 13 51 18
rect 21 11 51 13
rect 57 11 59 18
rect 69 16 71 18
rect 78 16 80 18
<< polycontact >>
rect 19 61 24 66
rect 27 57 31 61
rect 64 58 68 62
rect 32 30 37 35
rect 69 30 74 35
rect 12 6 16 11
rect 56 6 60 11
<< metal1 >>
rect -26 68 3 72
rect 7 68 17 72
rect 21 68 29 72
rect 35 68 53 72
rect 57 68 67 72
rect 72 68 81 72
rect 85 68 90 72
rect -26 66 90 68
rect 15 58 27 61
rect 15 54 19 58
rect 31 58 32 61
rect 16 53 19 54
rect 36 53 40 66
rect 51 58 64 61
rect 68 58 69 61
rect 51 54 55 58
rect 16 52 20 53
rect -20 44 -16 47
rect 0 44 4 47
rect 16 43 20 48
rect -20 24 -16 39
rect 0 24 4 39
rect 16 25 20 39
rect 25 47 29 48
rect 25 23 29 41
rect 52 53 55 54
rect 73 53 77 66
rect 52 52 56 53
rect 36 44 40 49
rect 44 43 48 48
rect 44 35 48 39
rect 37 30 48 35
rect 44 25 48 30
rect 52 43 56 48
rect 52 25 56 39
rect 62 47 66 48
rect 62 23 66 41
rect 73 44 77 49
rect 81 43 85 48
rect 81 35 85 39
rect 74 30 85 35
rect 81 25 85 30
rect 36 6 40 18
rect 73 6 77 18
rect -26 4 90 6
rect -26 0 1 4
rect 5 0 17 4
rect 21 0 36 4
rect 40 0 57 4
rect 61 0 79 4
rect 83 0 90 4
<< metal2 >>
rect -10 34 -6 52
rect 8 34 12 52
rect -10 30 12 34
rect -10 19 -6 30
rect 8 19 12 30
rect 19 11 24 66
rect 12 6 60 11
<< labels >>
rlabel metal1 14 70 14 70 5 vdd
rlabel polysilicon 14 55 14 55 1 clk_b
rlabel metal1 32 3 32 3 1 Gnd
rlabel polycontact 71 32 71 32 1 Q
rlabel polycontact 34 32 34 32 1 Q_b
rlabel metal2 14 8 14 8 1 clk
rlabel polysilicon -13 15 -13 15 1 s
rlabel polysilicon -14 62 -14 62 1 s_b
rlabel metal1 -18 33 -18 33 1 D
rlabel metal1 2 27 2 27 1 si
<< end >>
