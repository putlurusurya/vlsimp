magic
tech min2
timestamp 1606886706
<< error_p >>
rect -15 -7 -14 -3
rect -11 -7 -10 -3
<< nwell >>
rect -28 24 25 68
<< ntransistor >>
rect -13 1 -11 6
rect -8 1 -6 6
rect 1 1 3 6
rect 10 1 12 6
<< ptransistor >>
rect -13 47 -11 57
rect -8 47 -6 57
rect 1 47 3 57
rect 10 47 12 57
<< ndiffusion >>
rect -15 2 -13 6
rect -19 1 -13 2
rect -11 1 -8 6
rect -6 5 1 6
rect -6 1 -4 5
rect 0 1 1 5
rect 3 2 4 6
rect 9 2 10 6
rect 3 1 10 2
rect 12 5 18 6
rect 12 1 14 5
<< pdiffusion >>
rect -19 56 -13 57
rect -15 52 -13 56
rect -19 51 -13 52
rect -15 47 -13 51
rect -11 47 -8 57
rect -6 53 -4 57
rect 0 53 1 57
rect -6 52 1 53
rect -6 48 -4 52
rect 0 48 1 52
rect -6 47 1 48
rect 3 47 10 57
rect 12 56 18 57
rect 12 52 14 56
rect 12 51 18 52
rect 12 47 14 51
<< ndcontact >>
rect -19 2 -15 6
rect -4 1 0 5
rect 4 2 9 6
rect 14 1 18 5
<< pdcontact >>
rect -19 52 -15 56
rect -19 47 -15 51
rect -4 53 0 57
rect -4 48 0 52
rect 14 52 18 56
rect 14 47 18 51
<< psubstratepdiff >>
rect -11 -7 -7 -3
<< psubstratepcontact >>
rect -18 -7 -14 -3
rect 5 -7 9 -3
<< nsubstratencontact >>
rect -24 61 -20 65
rect -5 61 -1 65
rect 5 61 9 65
<< polysilicon >>
rect -13 57 -11 59
rect -8 57 -6 59
rect 1 57 3 59
rect 10 57 12 59
rect -13 45 -11 47
rect -8 45 -6 47
rect -13 41 -6 45
rect -13 12 -11 41
rect -8 31 -6 41
rect 1 39 3 47
rect 10 39 12 47
rect 2 35 3 39
rect 11 35 12 39
rect -8 27 -7 31
rect -8 12 -6 27
rect -13 8 -6 12
rect -13 6 -11 8
rect -8 6 -6 8
rect 1 6 3 35
rect 10 6 12 35
rect -13 -1 -11 1
rect -8 -1 -6 1
rect 1 -1 3 1
rect 10 -1 12 1
<< polycontact >>
rect -3 35 2 39
rect 6 35 11 39
rect -7 27 -2 31
<< metal1 >>
rect -25 61 -24 65
rect -20 61 -5 65
rect -1 61 5 65
rect 9 61 21 65
rect -25 59 21 61
rect -4 57 0 59
rect -19 51 -15 52
rect -4 52 0 53
rect 14 51 18 52
rect -19 28 -15 47
rect 14 31 18 47
rect -25 24 -15 28
rect -2 27 18 31
rect -19 6 -15 24
rect 5 6 8 27
rect -4 -1 0 1
rect 14 -1 18 1
rect -24 -3 21 -1
rect -24 -7 -18 -3
rect -14 -7 5 -3
rect 9 -7 21 -3
<< labels >>
rlabel metal1 2 -4 2 -4 1 Gnd
rlabel metal1 2 63 2 63 5 vdd
rlabel polycontact 8 37 8 37 1 b
rlabel metal1 -25 24 -25 28 3 out
rlabel polycontact 0 37 0 37 1 a
<< end >>
