magic
tech min2
timestamp 1606749416
<< nwell >>
rect -1 -12 153 33
<< ntransistor >>
rect 10 -26 12 -21
rect 30 -26 32 -21
rect 38 -26 40 -21
rect 46 -26 48 -21
rect 55 -26 57 -21
rect 63 -26 65 -21
rect 71 -26 73 -21
rect 101 -26 103 -21
rect 128 -26 130 -21
rect 136 -26 138 -21
<< ptransistor >>
rect 10 -1 12 9
rect 30 -1 32 9
rect 38 -1 40 9
rect 46 -1 48 9
rect 55 -1 57 9
rect 63 -1 65 9
rect 71 -1 73 9
rect 101 -1 103 9
rect 128 -6 130 12
rect 136 -6 138 12
<< ndiffusion >>
rect 5 -22 10 -21
rect 9 -26 10 -22
rect 12 -25 13 -21
rect 12 -26 17 -25
rect 29 -25 30 -21
rect 25 -26 30 -25
rect 32 -25 33 -21
rect 37 -25 38 -21
rect 32 -26 38 -25
rect 40 -25 41 -21
rect 45 -25 46 -21
rect 40 -26 46 -25
rect 48 -22 55 -21
rect 48 -26 50 -22
rect 54 -26 55 -22
rect 57 -25 58 -21
rect 62 -25 63 -21
rect 57 -26 63 -25
rect 65 -25 66 -21
rect 70 -25 71 -21
rect 65 -26 71 -25
rect 73 -25 74 -21
rect 73 -26 78 -25
rect 100 -25 101 -21
rect 96 -26 101 -25
rect 103 -22 108 -21
rect 103 -26 104 -22
rect 123 -22 128 -21
rect 127 -26 128 -22
rect 130 -25 131 -21
rect 135 -25 136 -21
rect 130 -26 136 -25
rect 138 -22 143 -21
rect 138 -26 139 -22
<< pdiffusion >>
rect 5 4 10 9
rect 9 0 10 4
rect 5 -1 10 0
rect 12 8 17 9
rect 12 4 13 8
rect 12 -1 17 4
rect 25 8 30 9
rect 29 4 30 8
rect 25 -1 30 4
rect 32 8 38 9
rect 32 4 33 8
rect 37 4 38 8
rect 32 -1 38 4
rect 40 8 46 9
rect 40 4 41 8
rect 45 4 46 8
rect 40 -1 46 4
rect 48 4 55 9
rect 48 0 50 4
rect 54 0 55 4
rect 48 -1 55 0
rect 57 8 63 9
rect 57 4 58 8
rect 62 4 63 8
rect 57 -1 63 4
rect 65 8 71 9
rect 65 4 66 8
rect 70 4 71 8
rect 65 -1 71 4
rect 73 8 78 9
rect 73 4 74 8
rect 73 -1 78 4
rect 96 8 101 9
rect 100 4 101 8
rect 96 -1 101 4
rect 103 4 108 9
rect 103 0 104 4
rect 103 -1 108 0
rect 123 8 128 12
rect 127 4 128 8
rect 123 3 128 4
rect 127 -1 128 3
rect 123 -6 128 -1
rect 130 -6 136 12
rect 138 9 143 12
rect 138 5 139 9
rect 138 4 143 5
rect 138 0 139 4
rect 138 -6 143 0
<< ndcontact >>
rect 5 -26 9 -22
rect 13 -25 17 -21
rect 25 -25 29 -21
rect 33 -25 37 -21
rect 41 -25 45 -21
rect 50 -26 54 -22
rect 58 -25 62 -21
rect 66 -25 70 -21
rect 74 -25 78 -21
rect 96 -25 100 -21
rect 104 -26 108 -22
rect 123 -26 127 -22
rect 131 -25 135 -21
rect 139 -26 143 -22
<< pdcontact >>
rect 5 0 9 4
rect 13 4 17 8
rect 25 4 29 8
rect 33 4 37 8
rect 41 4 45 8
rect 50 0 54 4
rect 58 4 62 8
rect 66 4 70 8
rect 74 4 78 8
rect 96 4 100 8
rect 104 0 108 4
rect 123 4 127 8
rect 123 -1 127 3
rect 139 5 143 9
rect 139 0 143 4
<< psubstratepcontact >>
rect 4 -43 8 -39
rect 16 -43 20 -39
rect 30 -43 34 -39
rect 45 -43 49 -39
rect 60 -43 64 -39
rect 76 -43 80 -39
rect 94 -43 98 -39
rect 111 -43 115 -39
rect 127 -43 131 -39
rect 139 -43 143 -39
<< nsubstratencontact >>
rect 8 25 12 29
rect 25 25 29 29
rect 45 25 49 29
rect 63 25 67 29
rect 77 25 81 29
rect 95 25 99 29
rect 112 25 116 29
rect 129 25 133 29
<< polysilicon >>
rect 38 21 65 23
rect 10 16 32 18
rect 10 9 12 16
rect 30 9 32 16
rect 38 9 40 21
rect 47 15 57 18
rect 46 9 48 11
rect 55 9 57 15
rect 63 9 65 21
rect 96 15 130 18
rect 71 12 83 14
rect 128 12 130 15
rect 136 12 138 14
rect 71 9 73 12
rect 10 -21 12 -1
rect 30 -3 32 -1
rect 10 -34 12 -26
rect 19 -29 21 -6
rect 38 -10 40 -1
rect 30 -12 40 -10
rect 30 -21 32 -12
rect 38 -21 40 -19
rect 46 -21 48 -1
rect 55 -21 57 -1
rect 63 -7 65 -1
rect 71 -3 73 -1
rect 63 -9 73 -7
rect 63 -21 65 -19
rect 71 -21 73 -9
rect 30 -29 32 -26
rect 19 -31 32 -29
rect 38 -34 40 -26
rect 46 -29 48 -26
rect 55 -29 57 -26
rect 63 -34 65 -26
rect 71 -29 73 -26
rect 81 -34 83 12
rect 101 9 103 11
rect 101 -21 103 -1
rect 128 -21 130 -6
rect 136 -9 138 -6
rect 136 -12 141 -9
rect 136 -21 138 -12
rect 101 -29 103 -26
rect 128 -29 130 -26
rect 136 -29 138 -26
rect 10 -36 83 -34
<< polycontact >>
rect 43 14 47 18
rect 92 15 96 19
rect 6 -18 10 -14
rect 15 -10 19 -6
rect 48 -12 52 -8
rect 103 -12 107 -8
rect 141 -12 146 -8
<< metal1 >>
rect 2 25 8 29
rect 12 25 25 29
rect 29 25 45 29
rect 49 25 63 29
rect 67 25 77 29
rect 81 25 95 29
rect 99 25 112 29
rect 116 25 129 29
rect 133 25 150 29
rect 2 23 150 25
rect 5 4 9 23
rect 33 15 43 18
rect 33 8 37 15
rect 13 -6 17 4
rect 13 -10 15 -6
rect 25 -8 29 4
rect 5 -18 6 -14
rect 13 -21 17 -10
rect 24 -12 29 -8
rect 25 -21 29 -12
rect 33 -21 37 4
rect 41 -21 45 4
rect 50 4 54 23
rect 58 15 92 18
rect 58 8 62 15
rect 58 -9 62 4
rect 52 -12 62 -9
rect 58 -21 62 -12
rect 5 -37 9 -26
rect 66 -21 70 4
rect 74 -9 78 4
rect 88 -9 91 -5
rect 96 -9 100 4
rect 104 4 108 23
rect 139 9 143 23
rect 123 3 127 4
rect 139 4 143 5
rect 74 -12 100 -9
rect 114 -9 117 -5
rect 123 -9 127 -1
rect 107 -12 135 -9
rect 146 -12 150 -9
rect 74 -21 78 -12
rect 96 -21 100 -12
rect 131 -21 135 -12
rect 50 -37 54 -26
rect 104 -37 108 -26
rect 123 -37 127 -26
rect 139 -37 143 -26
rect 2 -39 150 -37
rect 2 -43 4 -39
rect 8 -43 16 -39
rect 20 -43 30 -39
rect 34 -43 45 -39
rect 49 -43 60 -39
rect 64 -43 76 -39
rect 80 -43 94 -39
rect 98 -43 111 -39
rect 115 -43 127 -39
rect 131 -43 139 -39
rect 143 -43 150 -39
<< labels >>
rlabel polycontact 8 -16 8 -16 1 clk
rlabel metal1 25 -10 25 -10 1 D
rlabel metal1 115 -7 115 -7 1 Q
rlabel metal1 90 -7 90 -7 1 QB
rlabel pdcontact 7 2 7 2 3 t1
rlabel pdcontact 15 6 15 6 1 t2
rlabel pdcontact 27 6 27 6 1 t7
rlabel pdcontact 35 6 35 6 1 t8
rlabel pdcontact 43 6 43 6 1 t9
rlabel pdcontact 52 2 52 2 1 t10
rlabel pdcontact 60 6 60 6 1 t13
rlabel pdcontact 68 6 68 6 1 t14
rlabel pdcontact 76 6 76 6 1 t18
rlabel pdcontact 98 6 98 6 1 t21
rlabel pdcontact 106 2 106 2 1 t22
rlabel pdcontact 125 6 125 6 1 t23
rlabel pdcontact 142 2 142 2 1 t26
rlabel polycontact 144 -10 144 -10 1 clr
rlabel metal1 73 26 73 26 5 vdd
rlabel metal1 73 -41 73 -41 1 Gnd
rlabel ndcontact 7 -24 7 -24 3 t3
rlabel ndcontact 15 -23 15 -23 1 t4
rlabel ndcontact 27 -23 27 -23 1 t5
rlabel ndcontact 35 -23 35 -23 1 t6
rlabel ndcontact 43 -23 43 -23 1 t11
rlabel ndcontact 52 -24 52 -24 1 t12
rlabel ndcontact 60 -23 60 -23 1 t15
rlabel ndcontact 68 -23 68 -23 1 t16
rlabel ndcontact 76 -23 76 -23 1 t17
rlabel ndcontact 98 -23 98 -23 1 t19
rlabel ndcontact 107 -24 107 -24 1 t20
rlabel ndcontact 125 -24 125 -24 1 t24
rlabel ndcontact 133 -23 133 -23 1 t25
rlabel ndcontact 141 -24 141 -24 1 t24
<< end >>
