magic
tech min2
timestamp 1606882456
<< nwell >>
rect -44 24 28 69
<< ntransistor >>
rect -24 1 -22 6
rect -6 1 -4 6
rect 2 1 4 6
rect 11 1 13 6
<< ptransistor >>
rect -24 47 -22 57
rect -6 47 -4 57
rect 2 47 4 57
rect 11 47 13 57
<< ndiffusion >>
rect -26 2 -24 6
rect -30 1 -24 2
rect -22 5 -16 6
rect -22 1 -20 5
rect -8 2 -6 6
rect -12 1 -6 2
rect -4 5 2 6
rect -4 1 -3 5
rect 1 1 2 5
rect 4 1 11 6
rect 13 2 14 6
rect 13 1 18 2
<< pdiffusion >>
rect -30 56 -24 57
rect -26 52 -24 56
rect -30 51 -24 52
rect -26 47 -24 51
rect -22 53 -20 57
rect -22 52 -16 53
rect -22 48 -20 52
rect -22 47 -16 48
rect -12 56 -6 57
rect -8 52 -6 56
rect -12 51 -6 52
rect -8 47 -6 51
rect -4 52 2 57
rect -4 48 -3 52
rect 1 48 2 52
rect -4 47 2 48
rect 4 55 11 57
rect 4 51 5 55
rect 10 51 11 55
rect 4 47 11 51
rect 13 52 18 57
rect 13 48 14 52
rect 13 47 18 48
<< ndcontact >>
rect -30 2 -26 6
rect -20 1 -16 5
rect -12 2 -8 6
rect -3 1 1 5
rect 14 2 18 6
<< pdcontact >>
rect -30 52 -26 56
rect -30 47 -26 51
rect -20 53 -16 57
rect -20 48 -16 52
rect -12 52 -8 56
rect -12 47 -8 51
rect -3 48 1 52
rect 5 51 10 55
rect 14 48 18 52
<< psubstratepcontact >>
rect -41 -7 -37 -3
rect 6 -7 10 -3
rect 21 -7 25 -3
<< nsubstratencontact >>
rect -41 61 -37 65
rect 6 61 10 65
rect 21 61 25 65
<< polysilicon >>
rect -24 57 -22 59
rect -6 57 -4 59
rect 2 57 4 59
rect 11 57 13 59
rect -24 28 -22 47
rect -6 31 -4 47
rect -24 24 -23 28
rect -6 27 -5 31
rect -24 6 -22 24
rect -6 6 -4 27
rect 2 20 4 47
rect 3 16 4 20
rect 2 6 4 16
rect 11 6 13 47
rect -24 -1 -22 1
rect -6 -1 -4 1
rect 2 -1 4 1
rect 11 -1 13 1
<< polycontact >>
rect -23 24 -19 28
rect -5 27 -1 31
rect -1 16 3 20
rect 7 12 11 16
<< metal1 >>
rect -37 61 6 65
rect 10 61 21 65
rect -41 59 25 61
rect -20 57 -16 59
rect -30 51 -26 52
rect -20 52 -16 53
rect -12 51 -8 52
rect -30 28 -26 47
rect -3 52 1 59
rect 6 55 9 56
rect 14 52 18 59
rect -12 28 -8 47
rect 6 31 9 51
rect -33 24 -26 28
rect -19 24 -8 28
rect -1 27 18 31
rect -30 6 -26 24
rect -12 6 -8 24
rect -2 16 -1 20
rect 6 12 7 16
rect 14 6 18 27
rect -20 -1 -16 1
rect -3 -1 1 1
rect -41 -3 25 -1
rect -37 -7 6 -3
rect 10 -7 21 -3
<< labels >>
rlabel polycontact 9 14 9 14 1 b
rlabel metal1 3 -4 3 -4 1 Gnd
rlabel metal1 3 63 3 63 5 vdd
rlabel polycontact 1 18 1 18 1 a
rlabel metal1 -31 26 -31 26 1 out
<< end >>
