* SPICE3 file created from nor.ext - technology: min2

.option scale=0.1u

M1000 a_3_47# a vdd vdd pfet w=10 l=2
+  ad=70 pd=34 as=50 ps=30
M1001 out b a_3_47# vdd pfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1002 out a Gnd Gnd nfet w=5 l=2
+  ad=35 pd=24 as=50 ps=40
M1003 Gnd b out Gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
C0 out vdd 0.15456fF
C1 a vdd 0.23684fF
C2 a b 0.16295fF
C3 b vdd 0.23684fF


.include NMOS-180nm.lib
.include PMOS-180nm.lib


v_dd vdd Gnd 1.8
v_d a Gnd pulse( 1.8 0 0 1ns 1ns 50ns 100ns)

v1 b Gnd pulse(1.8 0 0 1ns 1ns 100ns 200ns)

.control
	tran 0.1ns 200ns
	
	plot tran1.a tran1.b tran1.out
	
	meas tran risetime  trig out val=0.18 RISE=1 TARG out val=1.62 RISE=1

	meas tran falltime  trig out val=1.62  FALL=1 TARG out val=0.18 FALL=1
	
	meas tran tplh trig a val=0.9 FALL=1 TARG out val=0.9 RISE=1
	
	meas tran tphl trig a val=0.9 RISE=1 TARG out val=0.9 FALL=1
	
	let x= -tran1.v_dd#branch
        
        plot vdd*x	   
	    
.endc

