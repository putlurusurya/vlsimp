* SPICE3 file created from nor.ext - technology: min2

.option scale=0.1u

M1000 a_n38_47# a_n40_n1# out vdd pfet w=10 l=2
+  ad=30 pd=26 as=50 ps=30
M1001 a_n33_47# a_n40_n1# a_n38_47# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1002 a_n28_47# a_n40_n1# a_n33_47# vdd pfet w=10 l=2
+  ad=30 pd=26 as=0 ps=0
M1003 vdd a_n40_n1# a_n28_47# vdd pfet w=10 l=2
+  ad=120 pd=64 as=0 ps=0
M1004 vdd a_n8_n1# a_n40_n1# vdd pfet w=10 l=2
+  ad=0 pd=0 as=60 ps=32
M1005 a_3_47# a vdd vdd pfet w=10 l=2
+  ad=70 pd=34 as=0 ps=0
M1006 a_n8_n1# b a_3_47# vdd pfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1007 a_n38_1# a_n40_n1# out Gnd nfet w=5 l=2
+  ad=15 pd=16 as=25 ps=20
M1008 a_n33_1# a_n40_n1# a_n38_1# Gnd nfet w=5 l=2
+  ad=15 pd=16 as=0 ps=0
M1009 a_n28_1# a_n40_n1# a_n33_1# Gnd nfet w=5 l=2
+  ad=15 pd=16 as=0 ps=0
M1010 Gnd a_n40_n1# a_n28_1# Gnd nfet w=5 l=2
+  ad=85 pd=64 as=0 ps=0
M1011 Gnd a_n8_n1# a_n40_n1# Gnd nfet w=5 l=2
+  ad=0 pd=0 as=30 ps=22
M1012 a_n8_n1# a Gnd Gnd nfet w=5 l=2
+  ad=35 pd=24 as=0 ps=0
M1013 Gnd b a_n8_n1# Gnd nfet w=5 l=2
+  ad=0 pd=0 as=0 ps=0
C0 b a 0.16295fF
C1 b a_n8_n1# 0.00719fF
C2 out vdd 0.16012fF
C3 a a_n8_n1# 0.18954fF
C4 a a_n40_n1# 0.02749fF
C5 b vdd 0.23684fF
C6 a_n8_n1# a_n40_n1# 0.05498fF
C7 a vdd 0.23684fF
C8 a_n8_n1# vdd 0.33938fF
C9 a_n40_n1# vdd 1.09350fF
C10 vdd Gnd 0.00263fF

.include NMOS-180nm.lib
.include PMOS-180nm.lib


v_dd vdd Gnd 1.8
v_d a Gnd pulse( 1.8 0 0 1ns 1ns 50ns 100ns)

v1 b Gnd pulse(1.8 0 0 1ns 1ns 100ns 200ns)

.control
	tran 0.1ns 200ns
	
	plot tran1.a tran1.b tran1.out
	
	meas tran risetime  trig out val=0.18 RISE=1 TARG out val=1.62 RISE=1

	meas tran falltime  trig out val=1.62  FALL=1 TARG out val=0.18 FALL=1
	
	meas tran tplh trig a val=0.9 FALL=1 TARG out val=0.9 RISE=1
	
	meas tran tphl trig a val=0.9 RISE=1 TARG out val=0.9 FALL=1
	
	let x= -tran1.v_dd#branch
        
        plot vdd*x	   
	    
.endc

