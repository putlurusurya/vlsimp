magic
tech min2
timestamp 1606885548
<< nwell >>
rect -23 24 26 69
<< ntransistor >>
rect -12 1 -10 6
rect -3 1 -1 6
rect 6 1 8 6
rect 11 1 13 6
<< ptransistor >>
rect -12 47 -10 57
rect -3 47 -1 57
rect 6 47 8 57
rect 11 47 13 57
<< ndiffusion >>
rect -13 2 -12 6
rect -17 1 -12 2
rect -10 1 -3 6
rect -1 5 6 6
rect -1 1 0 5
rect 4 1 6 5
rect 8 1 11 6
rect 13 2 14 6
rect 13 1 18 2
<< pdiffusion >>
rect -17 52 -12 57
rect -13 48 -12 52
rect -17 47 -12 48
rect -10 55 -3 57
rect -10 51 -9 55
rect -4 51 -3 55
rect -10 47 -3 51
rect -1 52 6 57
rect -1 48 0 52
rect 4 48 6 52
rect -1 47 6 48
rect 8 47 11 57
rect 13 56 18 57
rect 13 52 14 56
rect 13 51 18 52
rect 13 47 14 51
<< ndcontact >>
rect -17 2 -13 6
rect 0 1 4 5
rect 14 2 18 6
<< pdcontact >>
rect -17 48 -13 52
rect -9 51 -4 55
rect 0 48 4 52
rect 14 52 18 56
rect 14 47 18 51
<< psubstratepdiff >>
rect 7 -7 13 -3
<< nsubstratendiff >>
rect 7 61 14 65
<< psubstratepcontact >>
rect -9 -7 -5 -3
<< nsubstratencontact >>
rect -9 61 -5 65
<< polysilicon >>
rect -12 57 -10 59
rect -3 57 -1 59
rect 6 57 8 59
rect 11 57 13 60
rect -12 16 -10 47
rect -3 20 -1 47
rect 6 45 8 47
rect 11 45 13 47
rect 6 41 13 45
rect -3 16 -2 20
rect 6 16 8 41
rect 11 16 13 41
rect -12 12 -11 16
rect -12 6 -10 12
rect -3 6 -1 16
rect 6 12 13 16
rect 6 6 8 12
rect 11 6 13 12
rect -12 -1 -10 1
rect -3 -1 -1 1
rect 6 -1 8 1
rect 11 -1 13 1
<< polycontact >>
rect 2 27 6 31
rect -2 16 3 20
rect -11 12 -6 16
<< metal1 >>
rect -19 61 -9 65
rect -5 61 18 65
rect -19 60 18 61
rect -19 59 14 60
rect -17 52 -13 59
rect -8 55 -5 56
rect 0 52 4 59
rect -8 31 -5 51
rect 14 51 18 52
rect -18 27 2 31
rect 14 28 18 47
rect -18 6 -14 27
rect 14 24 26 28
rect 14 6 18 24
rect 0 -1 4 1
rect -19 -3 19 -1
rect -19 -7 -9 -3
rect -5 -7 19 -3
<< labels >>
rlabel metal1 -2 -4 -2 -4 1 Gnd
rlabel metal1 -2 63 -2 63 5 vdd
rlabel polycontact -9 14 -9 14 1 b
rlabel polycontact 1 18 1 18 1 a
rlabel metal1 21 25 21 25 7 out
<< end >>
