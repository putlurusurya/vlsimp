magic
tech min2
timestamp 1606748995
<< nwell >>
rect -14 24 27 69
<< ntransistor >>
rect 1 1 3 6
rect 10 1 12 6
<< ptransistor >>
rect 1 47 3 57
rect 10 47 12 57
<< ndiffusion >>
rect -4 5 1 6
rect 0 1 1 5
rect 3 1 10 6
rect 12 2 13 6
rect 12 1 17 2
<< pdiffusion >>
rect -4 52 1 57
rect 0 48 1 52
rect -4 47 1 48
rect 3 55 10 57
rect 3 51 4 55
rect 9 51 10 55
rect 3 47 10 51
rect 12 52 17 57
rect 12 48 13 52
rect 12 47 17 48
<< ndcontact >>
rect -4 1 0 5
rect 13 2 17 6
<< pdcontact >>
rect -4 48 0 52
rect 4 51 9 55
rect 13 48 17 52
<< psubstratepcontact >>
rect -11 -7 -7 -3
rect 5 -7 9 -3
rect 20 -7 24 -3
<< nsubstratencontact >>
rect -11 61 -7 65
rect 5 61 9 65
rect 20 61 24 65
<< polysilicon >>
rect 1 57 3 59
rect 10 57 12 59
rect 1 6 3 47
rect 10 6 12 47
rect 1 -1 3 1
rect 10 -1 12 1
<< polycontact >>
rect -3 16 1 20
rect 6 12 10 16
<< metal1 >>
rect -7 61 5 65
rect 9 61 20 65
rect -11 59 24 61
rect -4 52 0 59
rect 5 55 8 56
rect 13 52 17 59
rect 5 31 8 51
rect 5 27 24 31
rect -4 16 -3 20
rect 5 12 6 16
rect 13 6 17 27
rect -4 -1 0 1
rect -11 -3 24 -1
rect -7 -7 5 -3
rect 9 -7 20 -3
<< labels >>
rlabel polycontact 8 14 8 14 1 b
rlabel polycontact -1 18 -1 18 1 a
rlabel metal1 2 -4 2 -4 1 Gnd
rlabel metal1 24 27 24 31 7 out
rlabel metal1 2 63 2 63 5 vdd
<< end >>
